module sky130_fd_sc_hvl__lsbufhv2lv_1 (
    X,
    A
);

    output X;
    input  A;

    assign X = A;

endmodule